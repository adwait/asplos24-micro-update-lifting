
    module cache_ctrl_tb();
        parameter PHASE_TIME = 10;
        parameter CLK_CYCLE_TIME = PHASE_TIME * 2;
        parameter IMEM_INTERVAL = 20;
        parameter SIM_CYCLE = 21; // 100000000;
        parameter SIM_TIME = SIM_CYCLE * PHASE_TIME * 2;

        reg [31:0] 			CLK_CYCLE;
        reg 				clk;
        reg 				reset;
        
        initial begin
            clk = 1;
            forever #PHASE_TIME clk = ~clk;
        end

        initial begin
            reset = 1;
            // #IMEM_INTERVAL reset = 1;
            #IMEM_INTERVAL 
            reset = 0;
            #IMEM_INTERVAL 
            reset = 1;
        end
        
        initial begin
            CLK_CYCLE = 32'h0;
        end
        
        always @(posedge clk) begin
            CLK_CYCLE <= CLK_CYCLE + 1;
        end

        initial begin
            $dumpfile("cache_ctrl_wave_pipeline.vcd");
            $dumpvars(0, cache_ctrl_tb);
        end

        initial begin
            #IMEM_INTERVAL;
            #SIM_TIME;
            $finish;
        end


        // CSR tasks
        task make_tlb_lookup (input [19:0] vpn, input [8:0] asid);
            tb_io_update_i = 0;
            tb_io_lu_vaddr_i = {vpn, 12'h000};
            tb_io_lu_asid_i = asid;
            // Update stuff
            tb_io_flush_i = 0;
            tb_io_asid_to_be_flushed_i = 0;
            tb_io_vaddr_to_be_flushed_i = 0;
        endtask
        task make_tlb_update (input [19:0] vpn, input [8:0] asid, input [31:0] entry_data);
            tb_io_update_i = {1'b1, 1'b0, vpn, asid, entry_data};
            tb_io_lu_vaddr_i = 0;
            tb_io_lu_asid_i = 0;
            // Do not update anything
            tb_io_flush_i = 0;
            tb_io_asid_to_be_flushed_i = 0;
            tb_io_vaddr_to_be_flushed_i = 0;
        endtask
        task make_tlb_flush(input [19:0] vpn, input [8:0] asid);
            tb_io_update_i = 0;
            tb_io_lu_vaddr_i = 0;
            tb_io_lu_asid_i = 0;
            // Flush
            tb_io_flush_i = 1;
            tb_io_asid_to_be_flushed_i = asid;
            tb_io_vaddr_to_be_flushed_i = {vpn, 12'h000};
        endtask

        // Parameters and I/O connections
localparam ariane_pkg_NrMaxRules = 16;
localparam [6433:0] ariane_pkg_ArianeDefaultConfig =   
    6434'b10000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
parameter [6433:0] ArianeCfg = ariane_pkg_ArianeDefaultConfig;
localparam [31:0] ariane_pkg_CONFIG_L1D_SIZE = 32768;
localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = $clog2(32'd32768 / 32'd8);
localparam cva6_config_pkg_CVA6ConfigXlen = 32;
localparam riscv_XLEN = cva6_config_pkg_CVA6ConfigXlen;
localparam riscv_PLEN = 34;
localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = riscv_PLEN - ariane_pkg_DCACHE_INDEX_WIDTH;
localparam cva6_config_pkg_CVA6ConfigDataUserEn = 0;
localparam cva6_config_pkg_CVA6ConfigDataUserWidth = cva6_config_pkg_CVA6ConfigXlen;
localparam ariane_pkg_DATA_USER_WIDTH = 1;
localparam [31:0] ariane_pkg_DCACHE_USER_WIDTH = ariane_pkg_DATA_USER_WIDTH;
localparam [31:0] ariane_pkg_DCACHE_LINE_WIDTH = 128;
localparam std_cache_pkg_DCACHE_BYTE_OFFSET = 4;

        wire port_io_flush_i;
        reg tb_io_flush_i;
        assign port_io_flush_i = tb_io_flush_i;
        wire port_io_bypass_i;
        reg tb_io_bypass_i;
        assign port_io_bypass_i = tb_io_bypass_i;
        wire port_io_busy_o;
        wire [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + riscv_XLEN) + ariane_pkg_DCACHE_USER_WIDTH) + 9:0] port_io_req_port_i;
        reg [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + riscv_XLEN) + ariane_pkg_DCACHE_USER_WIDTH) + 9:0] tb_io_req_port_i;
        assign port_io_req_port_i = tb_io_req_port_i;
        reg [34:0] port_io_req_port_o;
        reg [7:0] port_io_req_o;
        reg [ariane_pkg_DCACHE_INDEX_WIDTH - 1:0] port_io_addr_o;
        wire port_io_gnt_i;
        reg tb_io_gnt_i;
        assign port_io_gnt_i = tb_io_gnt_i;
        reg [(ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 1:0] port_io_data_o;
        reg [((((ariane_pkg_DCACHE_TAG_WIDTH + 7) / 8) + 16) + ariane_pkg_DCACHE_SET_ASSOC) - 1:0] port_io_be_o;
        wire [ariane_pkg_DCACHE_TAG_WIDTH - 1:0] port_io_tag_o;
        wire [((ariane_pkg_DCACHE_TAG_WIDTH + 129) >= 0 ? (ariane_pkg_DCACHE_SET_ASSOC * ((ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 2)) - 1 : (ariane_pkg_DCACHE_SET_ASSOC * (1 - ((ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 1))) + ((ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 0)):((ariane_pkg_DCACHE_TAG_WIDTH + 129) >= 0 ? 0 : (ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 1)] port_io_data_i;
        reg [((ariane_pkg_DCACHE_TAG_WIDTH + 129) >= 0 ? (ariane_pkg_DCACHE_SET_ASSOC * ((ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 2)) - 1 : (ariane_pkg_DCACHE_SET_ASSOC * (1 - ((ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 1))) + ((ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 0)):((ariane_pkg_DCACHE_TAG_WIDTH + 129) >= 0 ? 0 : (ariane_pkg_DCACHE_TAG_WIDTH + ariane_pkg_DCACHE_LINE_WIDTH) + 1)] tb_io_data_i;
        assign tb_io_data_i = port_io_data_i;
        reg port_io_we_o;
        wire [7:0] port_io_hit_way_i;
        reg [7:0] tb_io_hit_way_i;
        assign port_io_hit_way_i = tb_io_hit_way_i;
        reg [140:0] port_io_miss_req_o;
        wire port_io_miss_gnt_i;
        reg tb_io_miss_gnt_i;
        assign port_io_miss_gnt_i = tb_io_miss_gnt_i;
        wire port_io_active_serving_i;
        reg tb_io_active_serving_i;
        assign port_io_active_serving_i = tb_io_active_serving_i;
        wire [63:0] port_io_critical_word_i;
        reg [63:0] tb_io_critical_word_i;
        assign port_io_critical_word_i = tb_io_critical_word_i;
        wire port_io_critical_word_valid_i;
        reg tb_io_critical_word_valid_i;
        assign port_io_critical_word_valid_i = tb_io_critical_word_valid_i;
        wire port_io_bypass_gnt_i;
        reg tb_io_bypass_gnt_i;
        assign port_io_bypass_gnt_i = tb_io_bypass_gnt_i;
        wire port_io_bypass_valid_i;
        reg tb_io_bypass_valid_i;
        assign port_io_bypass_valid_i = tb_io_bypass_valid_i;
        wire [63:0] port_io_bypass_data_i;
        reg [63:0] tb_io_bypass_data_i;
        assign port_io_bypass_data_i = tb_io_bypass_data_i;
        reg [55:0] port_io_mshr_addr_o;
        wire port_io_mshr_addr_matches_i;
        reg tb_io_mshr_addr_matches_i;
        assign port_io_mshr_addr_matches_i = tb_io_mshr_addr_matches_i;
        wire port_io_mshr_index_matches_i;
        reg tb_io_mshr_index_matches_i;
        assign port_io_mshr_index_matches_i = tb_io_mshr_index_matches_i;

        cache_ctrl cache_ctrl_i (
            .clk_i(clk),
	        .rst_ni(reset),
	        .flush_i(port_io_flush_i),
	        .bypass_i(port_io_bypass_i),
	        .busy_o(port_io_busy_o),
	        .req_port_i(port_io_req_port_i),
	        .req_port_o(port_io_req_port_o),
	        .req_o(port_io_req_o),
	        .addr_o(port_io_addr_o),
	        .gnt_i(port_io_gnt_i),
	        .data_o(port_io_data_o),
	        .be_o(port_io_be_o),
	        .tag_o(port_io_tag_o),
	        .data_i(port_io_data_i),
	        .we_o(port_io_we_o),
	        .hit_way_i(port_io_hit_way_i),
	        .miss_req_o(port_io_miss_req_o),
	        .miss_gnt_i(port_io_miss_gnt_i),
	        .active_serving_i(port_io_active_serving_i),
	        .critical_word_i(port_io_critical_word_i),
	        .critical_word_valid_i(port_io_critical_word_valid_i),
	        .bypass_gnt_i(port_io_bypass_gnt_i),
	        .bypass_valid_i(port_io_bypass_valid_i),
	        .bypass_data_i(port_io_bypass_data_i),
	        .mshr_addr_o(port_io_mshr_addr_o),
	        .mshr_addr_matches_i(port_io_mshr_addr_matches_i),
	        .mshr_index_matches_i(port_io_mshr_index_matches_i)
        );

        initial begin
            // Setup CSR
            #IMEM_INTERVAL;
            #IMEM_INTERVAL;
            #IMEM_INTERVAL;
            make_tlb_update(20'd10, 9'd1, 32'hffffffff);
            // make_csr_write(32'h0000007f, 32'hffffffff, 0);
            #20;
            make_tlb_lookup(20'd10, 9'd1);
            #20
            // make_csr_write(32'h00007f7f, 32'h00000000, 1);
            make_tlb_flush(0, 0);
            #20;
            make_tlb_lookup(20'd10, 9'd1);
        end
    endmodule
