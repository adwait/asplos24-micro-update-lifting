
    module ptw_tb();
        parameter PHASE_TIME = 10;
        parameter CLK_CYCLE_TIME = PHASE_TIME * 2;
        parameter IMEM_INTERVAL = 20;
        parameter SIM_CYCLE = 21; // 100000000;
        parameter SIM_TIME = SIM_CYCLE * PHASE_TIME * 2;

        reg [31:0] 			CLK_CYCLE;
        reg 				clk;
        reg 				reset;
        
        initial begin
            clk = 1;
            forever #PHASE_TIME clk = ~clk;
        end

        initial begin
            reset = 1;
            // #IMEM_INTERVAL reset = 1;
            #IMEM_INTERVAL 
            reset = 0;
            #IMEM_INTERVAL 
            reset = 1;
        end
        
        initial begin
            CLK_CYCLE = 32'h0;
        end
        
        always @(posedge clk) begin
            CLK_CYCLE <= CLK_CYCLE + 1;
        end

        initial begin
            $dumpfile("ptw_wave_pipeline.vcd");
            $dumpvars(0, ptw_tb);
        end

        initial begin
            #IMEM_INTERVAL;
            #SIM_TIME;
            $finish;
        end


        // CSR tasks
        task make_tlb_lookup (input [19:0] vpn, input [8:0] asid);
            tb_io_update_i = 0;
            tb_io_lu_vaddr_i = {vpn, 12'h000};
            tb_io_lu_asid_i = asid;
            // Update stuff
            tb_io_flush_i = 0;
            tb_io_asid_to_be_flushed_i = 0;
            tb_io_vaddr_to_be_flushed_i = 0;
        endtask
        task make_tlb_update (input [19:0] vpn, input [8:0] asid, input [31:0] entry_data);
            tb_io_update_i = {1'b1, 1'b0, vpn, asid, entry_data};
            tb_io_lu_vaddr_i = 0;
            tb_io_lu_asid_i = 0;
            // Do not update anything
            tb_io_flush_i = 0;
            tb_io_asid_to_be_flushed_i = 0;
            tb_io_vaddr_to_be_flushed_i = 0;
        endtask
        task make_tlb_flush(input [19:0] vpn, input [8:0] asid);
            tb_io_update_i = 0;
            tb_io_lu_vaddr_i = 0;
            tb_io_lu_asid_i = 0;
            // Flush
            tb_io_flush_i = 1;
            tb_io_asid_to_be_flushed_i = asid;
            tb_io_vaddr_to_be_flushed_i = {vpn, 12'h000};
        endtask

        // Parameters and I/O connections
localparam ariane_pkg_NrMaxRules = 16;
localparam [6433:0] ariane_pkg_ArianeDefaultConfig = 
    6434'b10000000000000000000000000001000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
localparam cva6_config_pkg_CVA6ConfigDataUserEn = 0;
localparam cva6_config_pkg_CVA6ConfigXlen = 32;
localparam cva6_config_pkg_CVA6ConfigDataUserWidth = cva6_config_pkg_CVA6ConfigXlen;
localparam ariane_pkg_DATA_USER_WIDTH = 1;
localparam [31:0] ariane_pkg_DCACHE_USER_WIDTH = ariane_pkg_DATA_USER_WIDTH;
localparam riscv_XLEN = cva6_config_pkg_CVA6ConfigXlen;
localparam [31:0] ariane_pkg_CONFIG_L1D_SIZE = 32768;
localparam [31:0] ariane_pkg_DCACHE_SET_ASSOC = 8;
localparam [31:0] ariane_pkg_DCACHE_INDEX_WIDTH = $clog2(32'd32768 / 32'd8);
localparam riscv_PLEN = 34;
localparam [31:0] ariane_pkg_DCACHE_TAG_WIDTH = riscv_PLEN - ariane_pkg_DCACHE_INDEX_WIDTH;
localparam riscv_VLEN = 32;
localparam riscv_PPNW = 22;
localparam [3:0] riscv_MODE_SV = 4'd1;
localparam riscv_SV = (riscv_MODE_SV == 4'd1 ? 32 : 39);
    
    // Flush the next instruction
    wire flush_i;
    reg tb_io_flush_i;
    assign port_io_flush_i = tb_io_flush_i;
    wire ptw_active_o;
    wire walking_instr_o;
    reg ptw_error_o;
    reg ptw_access_exception_o;
    
    // Disable address translation for instructions
    wire enable_translation_i;
    // reg tb_io_enable_translation_i;
    assign port_io_enable_translation_i = 0; // tb_io_enable_translation_i;
    // Always enable translation for loads and stores
    wire en_ld_st_translation_i;
    reg tb_io_en_ld_st_translation_i;
    assign port_io_en_ld_st_translation_i = 1; // tb_io_en_ld_st_translation_i;
    
    wire lsu_is_store_i;
    reg tb_io_lsu_is_store_i;
    assign port_io_lsu_is_store_i = tb_io_lsu_is_store_i;
    wire [34:0] req_port_i;
    reg [34:0] tb_io_req_port_i;
    assign port_io_req_port_i = tb_io_req_port_i;
    reg [(((ariane_pkg_DCACHE_INDEX_WIDTH + ariane_pkg_DCACHE_TAG_WIDTH) + riscv_XLEN) + ariane_pkg_DCACHE_USER_WIDTH) + 9:0] port_io_req_port_o;
    reg [62:0] itlb_update_o;
    reg [62:0] dtlb_update_o;
    wire [31:0] update_vaddr_o;
    wire [ASID_WIDTH - 1:0] asid_i;
    reg [ASID_WIDTH - 1:0] tb_io_asid_i;
    assign port_io_asid_i = tb_io_asid_i;
    
    // No accesses for instructions
    wire itlb_access_i;
    // reg tb_io_itlb_access_i;
    assign port_io_itlb_access_i = 0; // tb_io_itlb_access_i;
    wire itlb_hit_i;
    // reg tb_io_itlb_hit_i;
    assign port_io_itlb_hit_i = 0; // tb_io_itlb_hit_i;
    wire [31:0] itlb_vaddr_i;
    // reg [31:0] tb_io_itlb_vaddr_i;
    assign port_io_itlb_vaddr_i = 0; // tb_io_itlb_vaddr_i;
    
    // Following two lines indicate that the dtlb is being accessed
    wire dtlb_access_i;
    reg tb_io_dtlb_access_i;
    assign port_io_dtlb_access_i = tb_io_dtlb_access_i;
    wire dtlb_hit_i;
    reg tb_io_dtlb_hit_i;
    assign port_io_dtlb_hit_i = tb_io_dtlb_hit_i;
    
    // Following lines indicate the physsical page number and virtual address
    wire [31:0] dtlb_vaddr_i;
    reg [31:0] tb_io_dtlb_vaddr_i;
    assign port_io_dtlb_vaddr_i = tb_io_dtlb_vaddr_i;
    wire [21:0] satp_ppn_i;
    reg [21:0] tb_io_satp_ppn_i;
    assign port_io_satp_ppn_i = tb_io_satp_ppn_i;
    
    wire mxr_i;
    reg tb_io_mxr_i;
    assign port_io_mxr_i = tb_io_mxr_i;
    reg itlb_miss_o;
    reg dtlb_miss_o;
    // wire [127:0] pmpcfg_i;
    // reg [127:0] tb_io_pmpcfg_i;
    // assign port_io_pmpcfg_i = tb_io_pmpcfg_i;
    // wire [511:0] pmpaddr_i;
    // reg [511:0] tb_io_pmpaddr_i;
    // assign port_io_pmpaddr_i = tb_io_pmpaddr_i;
    wire [33:0] bad_paddr_o;

        cva6_ptw_sv32 ptw_i (
            .clk_i(clk),
            .rst_ni(reset),
            .flush_i(port_io_flush_i),
            .ptw_active_o(port_io_ptw_active_o),
            .walking_instr_o(port_io_walking_instr_o),
            .ptw_error_o(port_io_ptw_error_o),
            .ptw_access_exception_o(port_io_ptw_access_exception_o),
            .enable_translation_i(port_io_enable_translation_i),
            .en_ld_st_translation_i(port_io_en_ld_st_translation_i),
            .lsu_is_store_i(port_io_lsu_is_store_i),
            .req_port_i(port_io_req_port_i),
            .req_port_o(port_io_req_port_o),
            .itlb_update_o(port_io_itlb_update_o),
            .dtlb_update_o(port_io_dtlb_update_o),
            .update_vaddr_o(port_io_update_vaddr_o),
            .asid_i(port_io_asid_i),
            .itlb_access_i(port_io_itlb_access_i),
            .itlb_hit_i(port_io_itlb_hit_i),
            .itlb_vaddr_i(port_io_itlb_vaddr_i),
            .dtlb_access_i(port_io_dtlb_access_i),
            .dtlb_hit_i(port_io_dtlb_hit_i),
            .dtlb_vaddr_i(port_io_dtlb_vaddr_i),
            .satp_ppn_i(port_io_satp_ppn_i),
            .mxr_i(port_io_mxr_i),
            .itlb_miss_o(port_io_itlb_miss_o),
            .dtlb_miss_o(port_io_dtlb_miss_o),
            .pmpcfg_i(port_io_conf_i),
            .pmpaddr_i(port_io_conf_addr_i),
            .bad_paddr_o(port_io_bad_paddr_o),
        );

        simple_csr_regfile csr_f (
            .clk_i(clk),
            .rst_ni(reset),
            .csr_wdata_i(port_io_csr_wdata_i),
            .csr_addr_i(port_io_csr_addr_i),
            .csr_op_i(port_io_csr_op_i),
            .pmpcfg_o(port_io_conf_i),
            .pmpaddr_o(port_io_conf_addr_i)
        );

        initial begin
            // Setup CSR
            #IMEM_INTERVAL;
            #IMEM_INTERVAL;
            #IMEM_INTERVAL;
            make_tlb_update(20'd10, 9'd1, 32'hffffffff);
            // make_csr_write(32'h0000007f, 32'hffffffff, 0);
            #20;
            make_tlb_lookup(20'd10, 9'd1);
            #20
            // make_csr_write(32'h00007f7f, 32'h00000000, 1);
            make_tlb_flush(0, 0);
            #20;
            make_tlb_lookup(20'd10, 9'd1);
        end
    endmodule
